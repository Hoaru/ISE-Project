//----------------------------------------------
//ѡ����ģ��
//----------------------------------------------
module mux2(A,B,Z,s); 
input[31:0] A,B; 
input s;
output[31:0] Z;
wire[31:0] Z;
assign Z = (s == 1)?A:B;
endmodule
